module add2 (output logic [1:0] out, )
